module ROM(
    output reg[28:0] DataROM,
    input wire[10:0] AddrROM
);
    reg[28:0] data [2047:0];
    initial begin
        data[0] = 29'h01f040ff;
        data[1] = 29'h01000001;
        data[2] = 29'h15000008;
        data[3] = 29'h0100c5e8;
        data[4] = 29'h15000007;
        data[5] = 29'h01000048;
        data[6] = 29'h15004000;
        data[7] = 29'h1600f000;
        data[8] = 29'h05ff0001;
        data[9] = 29'h1200001f;
        data[10] = 29'h01000069;
        data[11] = 29'h15004000;
        data[12] = 29'h1600f000;
        data[13] = 29'h05ff0001;
        data[14] = 29'h1200001f;
        data[15] = 29'h0100003a;
        data[16] = 29'h15004000;
        data[17] = 29'h1600f000;
        data[18] = 29'h05ff0001;
        data[19] = 29'h1200001f;
        data[20] = 29'h01000020;
        data[21] = 29'h15004000;
        data[22] = 29'h1600f000;
        data[23] = 29'h05ff0001;
        data[24] = 29'h1200001f;
        data[25] = 29'h01008702;
        data[26] = 29'h15004000;
        data[27] = 29'h1600f000;
        data[28] = 29'h05ff0001;
        data[29] = 29'h1200002a;
        data[30] = 29'h1200001e;
        data[31] = 29'h18004000;
        data[32] = 29'h0f000100;
        data[33] = 29'h15000006;
        data[34] = 29'h0b00feff;
        data[35] = 29'h15000006;
        data[36] = 29'h18000009;
        data[37] = 29'h0b000002;
        data[38] = 29'h12010028;
        data[39] = 29'h12000024;
        data[40] = 29'h03ff0001;
        data[41] = 29'h1700f000;
        data[42] = 29'h01000000;
        data[43] = 29'h01100000;
        data[44] = 29'h18204000;
        data[45] = 29'h01300000;
        data[46] = 29'h01400000;
        data[47] = 29'h08a04000;
        data[48] = 29'h0baa000f;
        data[49] = 29'h05aa0005;
        data[50] = 29'h12030036;
        data[51] = 29'h01a00003;
        data[52] = 29'h06aa4000;
        data[53] = 29'h0200a000;
        data[54] = 29'h03440004;
        data[55] = 29'h05a40010;
        data[56] = 29'h1203002f;
        data[57] = 29'h0ba1000f;
        data[58] = 29'h05aa0005;
        data[59] = 29'h1203003d;
        data[60] = 29'h03110003;
        data[61] = 29'h07a10001;
        data[62] = 29'h09b0000f;
        data[63] = 29'h0e1ab000;
        data[64] = 29'h07a00001;
        data[65] = 29'h09b2000f;
        data[66] = 29'h0e0ab000;
        data[67] = 29'h07220001;
        data[68] = 29'h03330001;
        data[69] = 29'h05a30010;
        data[70] = 29'h1203002e;
        data[71] = 29'h0b81000f;
        data[72] = 29'h1201004d;
        data[73] = 29'h03880130;
        data[74] = 29'h15080006;
        data[75] = 29'h0b88003f;
        data[76] = 29'h15080006;
        data[77] = 29'h0b90f000;
        data[78] = 29'h02a98000;
        data[79] = 29'h12010055;
        data[80] = 29'h0989000c;
        data[81] = 29'h03880130;
        data[82] = 29'h15080006;
        data[83] = 29'h0b88003f;
        data[84] = 29'h15080006;
        data[85] = 29'h0ba00f00;
        data[86] = 29'h028a9000;
        data[87] = 29'h1201005d;
        data[88] = 29'h098a0008;
        data[89] = 29'h03880130;
        data[90] = 29'h15080006;
        data[91] = 29'h0b88003f;
        data[92] = 29'h15080006;
        data[93] = 29'h0bb000f0;
        data[94] = 29'h02aba000;
        data[95] = 29'h12010065;
        data[96] = 29'h098b0004;
        data[97] = 29'h03880130;
        data[98] = 29'h15080006;
        data[99] = 29'h0b88003f;
        data[100] = 29'h15080006;
        data[101] = 29'h0b80000f;
        data[102] = 29'h03880130;
        data[103] = 29'h15080006;
        data[104] = 29'h0b88003f;
        data[105] = 29'h15080006;
        data[106] = 29'h15004000;
        data[107] = 29'h15014001;
        data[108] = 29'h03ff0001;
        data[109] = 29'h1700f000;
    end
    
    // Lecture synchrone ou asynchrone de la ROM
    always @(*) begin
        DataROM = data[AddrROM];
    end
endmodule
