module ROM(
    output reg[28:0] DataROM,
    input wire[7:0] AddrROM
);
    reg[28:0] data [255:0];
    initial begin      
        data[0] = 29'h01000001;
        data[1] = 29'h15000007;
        data[2] = 29'h0100c5e8;
        data[3] = 29'h15000006;
        data[4] = 29'h01000143;
        data[5] = 29'h15000005;
        data[6] = 29'h01000000;
        data[7] = 29'h15000005;
        data[8] = 29'h01000161;
        data[9] = 29'h15000005;
        data[10] = 29'h01000000;
        data[11] = 29'h15000005;
        data[12] = 29'h0100016c;
        data[13] = 29'h15000005;
        data[14] = 29'h01000000;
        data[15] = 29'h15000005;
        data[16] = 29'h01000163;
        data[17] = 29'h15000005;
        data[18] = 29'h01000000;
        data[19] = 29'h15000005;
        data[20] = 29'h01000120;
        data[21] = 29'h15000005;
        data[22] = 29'h01000000;
        data[23] = 29'h15000005;
        data[24] = 29'h01000152;
        data[25] = 29'h15000005;
        data[26] = 29'h01000000;
        data[27] = 29'h15000005;
        data[28] = 29'h01000165;
        data[29] = 29'h15000005;
        data[30] = 29'h01000000;
        data[31] = 29'h15000005;
        data[32] = 29'h01000173;
        data[33] = 29'h15000005;
        data[34] = 29'h01000000;
        data[35] = 29'h15000005;
        data[36] = 29'h01000120;
        data[37] = 29'h15000005;
        data[38] = 29'h01000000;
        data[39] = 29'h15000005;
        data[40] = 29'h01000153;
        data[41] = 29'h15000005;
        data[42] = 29'h01000000;
        data[43] = 29'h15000005;
        data[44] = 29'h01000165;
        data[45] = 29'h15000005;
        data[46] = 29'h01000000;
        data[47] = 29'h15000005;
        data[48] = 29'h01000172;
        data[49] = 29'h15000005;
        data[50] = 29'h01000000;
        data[51] = 29'h15000005;
        data[52] = 29'h01000169;
        data[53] = 29'h15000005;
        data[54] = 29'h01000000;
        data[55] = 29'h15000005;
        data[56] = 29'h01000165;
        data[57] = 29'h15000005;
        data[58] = 29'h01000000;
        data[59] = 29'h15000005;
        data[60] = 29'h0100013a;
        data[61] = 29'h15000005;
        data[62] = 29'h01000000;
        data[63] = 29'h15000005;
        data[64] = 29'h0100010a;
        data[65] = 29'h01100000;
        data[66] = 29'h15000005;
        data[67] = 29'h15010005;
        data[68] = 29'h0100010d;
        data[69] = 29'h15000005;
        data[70] = 29'h15010005;
        data[71] = 29'h0100010a;
        data[72] = 29'h01100000;
        data[73] = 29'h15000005;
        data[74] = 29'h15010005;
        data[75] = 29'h0100010d;
        data[76] = 29'h15000005;
        data[77] = 29'h15010005;
        data[78] = 29'h01000152;
        data[79] = 29'h15000005;
        data[80] = 29'h01000000;
        data[81] = 29'h15000005;
        data[82] = 29'h01000131;
        data[83] = 29'h15000005;
        data[84] = 29'h01000000;
        data[85] = 29'h15000005;
        data[86] = 29'h0100013a;
        data[87] = 29'h15000005;
        data[88] = 29'h01000000;
        data[89] = 29'h15000005;
        data[90] = 29'h01000120;
        data[91] = 29'h15000005;
        data[92] = 29'h01000000;
        data[93] = 29'h15000005;
        data[94] = 29'h01800000;
        data[95] = 29'h01000005;
        data[96] = 29'h13800000;
        data[97] = 29'h05780030;
        data[98] = 29'h1203005e;
        data[99] = 29'h03080100;
        data[100] = 29'h15000005;
        data[101] = 29'h01000000;
        data[102] = 29'h15000005;
        data[103] = 29'h0100010a;
        data[104] = 29'h01100000;
        data[105] = 29'h15000005;
        data[106] = 29'h15010005;
        data[107] = 29'h0100010d;
        data[108] = 29'h15000005;
        data[109] = 29'h15010005;
        data[110] = 29'h01000152;
        data[111] = 29'h15000005;
        data[112] = 29'h01000000;
        data[113] = 29'h15000005;
        data[114] = 29'h01000132;
        data[115] = 29'h15000005;
        data[116] = 29'h01000000;
        data[117] = 29'h15000005;
        data[118] = 29'h0100013a;
        data[119] = 29'h15000005;
        data[120] = 29'h01000000;
        data[121] = 29'h15000005;
        data[122] = 29'h01000120;
        data[123] = 29'h15000005;
        data[124] = 29'h01000000;
        data[125] = 29'h15000005;
        data[126] = 29'h01900000;
        data[127] = 29'h01000005;
        data[128] = 29'h13900000;
        data[129] = 29'h05790030;
        data[130] = 29'h1203007e;
        data[131] = 29'h03090100;
        data[132] = 29'h15000005;
        data[133] = 29'h01000000;
        data[134] = 29'h15000005;
        data[135] = 29'h0100010a;
        data[136] = 29'h01100000;
        data[137] = 29'h15000005;
        data[138] = 29'h15010005;
        data[139] = 29'h0100010d;
        data[140] = 29'h15000005;
        data[141] = 29'h15010005;
        data[142] = 29'h01000152;
        data[143] = 29'h15000005;
        data[144] = 29'h01000000;
        data[145] = 29'h15000005;
        data[146] = 29'h01000165;
        data[147] = 29'h15000005;
        data[148] = 29'h01000000;
        data[149] = 29'h15000005;
        data[150] = 29'h01000171;
        data[151] = 29'h15000005;
        data[152] = 29'h01000000;
        data[153] = 29'h15000005;
        data[154] = 29'h01000120;
        data[155] = 29'h15000005;
        data[156] = 29'h01000000;
        data[157] = 29'h15000005;
        data[158] = 29'h0100013a;
        data[159] = 29'h15000005;
        data[160] = 29'h01000000;
        data[161] = 29'h15000005;
        data[162] = 29'h05690030;
        data[163] = 29'h02786000;
        data[164] = 29'h05070030;
        data[165] = 29'h15000002;
        data[166] = 29'h03070100;
        data[167] = 29'h15000005;
        data[168] = 29'h01000000;
        data[169] = 29'h15000005;
        data[170] = 29'h0100010a;
        data[171] = 29'h01100000;
        data[172] = 29'h15000005;
        data[173] = 29'h15010005;
        data[174] = 29'h0100010d;
        data[175] = 29'h15000005;
        data[176] = 29'h15010005;
        data[177] = 29'h0500000a;
        data[178] = 29'h120300b6;
        data[179] = 29'h03000061;
        data[180] = 29'h120000b7;
        data[181] = 29'h0300003a;
        data[182] = 29'h03000100;
        data[183] = 29'h15000005;
        data[184] = 29'h01000000;
        data[185] = 29'h15000005;
        data[186] = 29'h00000000;
        data[187] = 29'h00000000;
        data[188] = 29'h00000000;
        data[189] = 29'h00000000;
        data[190] = 29'h00000000;
        data[191] = 29'h00000000;
        data[192] = 29'h00000000;
        data[193] = 29'h00000000;
        data[194] = 29'h00000000;
        data[195] = 29'h00000000;
        data[196] = 29'h00000000;
        data[197] = 29'h00000000;
        data[198] = 29'h00000000;
        data[199] = 29'h00000000;
        data[200] = 29'h00000000;
        data[201] = 29'h00000000;
        data[202] = 29'h00000000;
        data[203] = 29'h00000000;
        data[204] = 29'h00000000;
        data[205] = 29'h00000000;
        data[206] = 29'h00000000;
        data[207] = 29'h00000000;
        data[208] = 29'h00000000;
        data[209] = 29'h00000000;
        data[210] = 29'h00000000;
        data[211] = 29'h00000000;
        data[212] = 29'h00000000;
        data[213] = 29'h00000000;
        data[214] = 29'h00000000;
        data[215] = 29'h00000000;
        data[216] = 29'h00000000;
        data[217] = 29'h00000000;
        data[218] = 29'h00000000;
        data[219] = 29'h00000000;
        data[220] = 29'h00000000;
        data[221] = 29'h00000000;
        data[222] = 29'h00000000;
        data[223] = 29'h00000000;
        data[224] = 29'h00000000;
        data[225] = 29'h00000000;
        data[226] = 29'h00000000;
        data[227] = 29'h00000000;
        data[228] = 29'h00000000;
        data[229] = 29'h00000000;
        data[230] = 29'h00000000;
        data[231] = 29'h00000000;
        data[232] = 29'h00000000;
        data[233] = 29'h00000000;
        data[234] = 29'h00000000;
        data[235] = 29'h00000000;
        data[236] = 29'h00000000;
        data[237] = 29'h00000000;
        data[238] = 29'h00000000;
        data[239] = 29'h00000000;
        data[240] = 29'h00000000;
        data[241] = 29'h00000000;
        data[242] = 29'h00000000;
        data[243] = 29'h00000000;
        data[244] = 29'h00000000;
        data[245] = 29'h00000000;
        data[246] = 29'h00000000;
        data[247] = 29'h00000000;
        data[248] = 29'h12000000;
        data[249] = 29'h12000000;
        data[250] = 29'h12000000;
        data[251] = 29'h12000000;
        data[252] = 29'h12000000;
        data[253] = 29'h12000000;
        data[254] = 29'h12000000;
        data[255] = 29'h12000000;
    end
    
// Lecture synchrone ou asynchrone de la ROM
    always @(*) begin
        DataROM = data[AddrROM];
    end
endmodule
