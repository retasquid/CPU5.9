module ROM(
    output reg[28:0] DataROM,
    input wire[10:0] AddrROM
);
    reg[28:0] data [2047:0];
    initial begin
        data[0] = 29'h01f0c0ff;
        data[1] = 29'h01000000;
        data[2] = 29'h15000008;
        data[3] = 29'h01002580;
        data[4] = 29'h15000007;
        data[5] = 29'h010000aa;
        data[6] = 29'h15000002;
        data[7] = 29'h1600f002;
        data[8] = 29'h05ff0001;
        data[9] = 29'h12000125;
        data[10] = 29'h01108000;
        data[11] = 29'h01001fff;
        data[12] = 29'h14001000;
        data[13] = 29'h03110001;
        data[14] = 29'h05000001;
        data[15] = 29'h12010011;
        data[16] = 29'h1200000c;
        data[17] = 29'h14001000;
        data[18] = 29'h01708000;
        data[19] = 29'h13007000;
        data[20] = 29'h05800000;
        data[21] = 29'h12010023;
        data[22] = 29'h1600f002;
        data[23] = 29'h05ff0001;
        data[24] = 29'h120000ab;
        data[25] = 29'h03770010;
        data[26] = 29'h0100000d;
        data[27] = 29'h1600f002;
        data[28] = 29'h05ff0001;
        data[29] = 29'h12000091;
        data[30] = 29'h0100000a;
        data[31] = 29'h1600f002;
        data[32] = 29'h05ff0001;
        data[33] = 29'h12000091;
        data[34] = 29'h12000013;
        data[35] = 29'h01000046;
        data[36] = 29'h1600f002;
        data[37] = 29'h05ff0001;
        data[38] = 29'h12000091;
        data[39] = 29'h01000069;
        data[40] = 29'h1600f002;
        data[41] = 29'h05ff0001;
        data[42] = 29'h12000091;
        data[43] = 29'h0100006e;
        data[44] = 29'h1600f002;
        data[45] = 29'h05ff0001;
        data[46] = 29'h12000091;
        data[47] = 29'h01000020;
        data[48] = 29'h1600f002;
        data[49] = 29'h05ff0001;
        data[50] = 29'h12000091;
        data[51] = 29'h01000064;
        data[52] = 29'h1600f002;
        data[53] = 29'h05ff0001;
        data[54] = 29'h12000091;
        data[55] = 29'h01000075;
        data[56] = 29'h1600f002;
        data[57] = 29'h05ff0001;
        data[58] = 29'h12000091;
        data[59] = 29'h01000020;
        data[60] = 29'h1600f002;
        data[61] = 29'h05ff0001;
        data[62] = 29'h12000091;
        data[63] = 29'h01000074;
        data[64] = 29'h1600f002;
        data[65] = 29'h05ff0001;
        data[66] = 29'h12000091;
        data[67] = 29'h01000065;
        data[68] = 29'h1600f002;
        data[69] = 29'h05ff0001;
        data[70] = 29'h12000091;
        data[71] = 29'h01000073;
        data[72] = 29'h1600f002;
        data[73] = 29'h05ff0001;
        data[74] = 29'h12000091;
        data[75] = 29'h01000074;
        data[76] = 29'h1600f002;
        data[77] = 29'h05ff0001;
        data[78] = 29'h12000091;
        data[79] = 29'h0100002c;
        data[80] = 29'h1600f002;
        data[81] = 29'h05ff0001;
        data[82] = 29'h12000091;
        data[83] = 29'h01000020;
        data[84] = 29'h1600f002;
        data[85] = 29'h05ff0001;
        data[86] = 29'h12000091;
        data[87] = 29'h01000053;
        data[88] = 29'h1600f002;
        data[89] = 29'h05ff0001;
        data[90] = 29'h12000091;
        data[91] = 29'h01000055;
        data[92] = 29'h1600f002;
        data[93] = 29'h05ff0001;
        data[94] = 29'h12000091;
        data[95] = 29'h01000043;
        data[96] = 29'h1600f002;
        data[97] = 29'h05ff0001;
        data[98] = 29'h12000091;
        data[99] = 29'h01000043;
        data[100] = 29'h1600f002;
        data[101] = 29'h05ff0001;
        data[102] = 29'h12000091;
        data[103] = 29'h01000045;
        data[104] = 29'h1600f002;
        data[105] = 29'h05ff0001;
        data[106] = 29'h12000091;
        data[107] = 29'h01000053;
        data[108] = 29'h1600f002;
        data[109] = 29'h05ff0001;
        data[110] = 29'h12000091;
        data[111] = 29'h010000ff;
        data[112] = 29'h15000002;
        data[113] = 29'h01002710;
        data[114] = 29'h1600f002;
        data[115] = 29'h05ff0001;
        data[116] = 29'h12000120;
        data[117] = 29'h01000000;
        data[118] = 29'h15000002;
        data[119] = 29'h01002710;
        data[120] = 29'h1600f002;
        data[121] = 29'h05ff0001;
        data[122] = 29'h12000120;
        data[123] = 29'h1200006f;
        data[124] = 29'h0ab11000;
        data[125] = 29'h18000006;
        data[126] = 29'h05000000;
        data[127] = 29'h1201007c;
        data[128] = 29'h05a0000d;
        data[129] = 29'h1201008d;
        data[130] = 29'h05a00008;
        data[131] = 29'h12010087;
        data[132] = 29'h14001000;
        data[133] = 29'h03110001;
        data[134] = 29'h12000089;
        data[135] = 29'h05110001;
        data[136] = 29'h140a1000;
        data[137] = 29'h1600f002;
        data[138] = 29'h05ff0001;
        data[139] = 29'h12000091;
        data[140] = 29'h1200007c;
        data[141] = 29'h140a1000;
        data[142] = 29'h0a0bb000;
        data[143] = 29'h03ff0001;
        data[144] = 29'h1700f000;
        data[145] = 29'h0f000100;
        data[146] = 29'h15000006;
        data[147] = 29'h0b00feff;
        data[148] = 29'h15000006;
        data[149] = 29'h18000009;
        data[150] = 29'h0b000002;
        data[151] = 29'h12010099;
        data[152] = 29'h12000095;
        data[153] = 29'h03ff0001;
        data[154] = 29'h1700f000;
        data[155] = 29'h01a00000;
        data[156] = 29'h01b00000;
        data[157] = 29'h13c00000;
        data[158] = 29'h03000001;
        data[159] = 29'h05cc0000;
        data[160] = 29'h120100a8;
        data[161] = 29'h07da0003;
        data[162] = 29'h07ea0001;
        data[163] = 29'h02dde000;
        data[164] = 29'h05cc0030;
        data[165] = 29'h02adc000;
        data[166] = 29'h03bb0001;
        data[167] = 29'h1200009d;
        data[168] = 29'h0a0aa000;
        data[169] = 29'h03ff0001;
        data[170] = 29'h1700f000;
        data[171] = 29'h0a200000;
        data[172] = 29'h01000000;
        data[173] = 29'h01100000;
        data[174] = 29'h01300000;
        data[175] = 29'h01400000;
        data[176] = 29'h08a04000;
        data[177] = 29'h0baa000f;
        data[178] = 29'h05aa0005;
        data[179] = 29'h120300b7;
        data[180] = 29'h01a00003;
        data[181] = 29'h06aa4000;
        data[182] = 29'h0200a000;
        data[183] = 29'h03440004;
        data[184] = 29'h05a40010;
        data[185] = 29'h120300b0;
        data[186] = 29'h0ba1000f;
        data[187] = 29'h05aa0005;
        data[188] = 29'h120300be;
        data[189] = 29'h03110003;
        data[190] = 29'h07a10001;
        data[191] = 29'h09b0000f;
        data[192] = 29'h0e1ab000;
        data[193] = 29'h07a00001;
        data[194] = 29'h09b2000f;
        data[195] = 29'h0e0ab000;
        data[196] = 29'h07220001;
        data[197] = 29'h03330001;
        data[198] = 29'h05a30010;
        data[199] = 29'h120300af;
        data[200] = 29'h0b81000f;
        data[201] = 29'h120100cd;
        data[202] = 29'h1600f002;
        data[203] = 29'h05ff0001;
        data[204] = 29'h120000e8;
        data[205] = 29'h0b90f000;
        data[206] = 29'h02a98000;
        data[207] = 29'h120100d4;
        data[208] = 29'h0989000c;
        data[209] = 29'h1600f002;
        data[210] = 29'h05ff0001;
        data[211] = 29'h120000e8;
        data[212] = 29'h0b900f00;
        data[213] = 29'h02aa9000;
        data[214] = 29'h120100db;
        data[215] = 29'h09890008;
        data[216] = 29'h1600f002;
        data[217] = 29'h05ff0001;
        data[218] = 29'h120000e8;
        data[219] = 29'h0b9000f0;
        data[220] = 29'h02a9a000;
        data[221] = 29'h120100e2;
        data[222] = 29'h09890004;
        data[223] = 29'h1600f002;
        data[224] = 29'h05ff0001;
        data[225] = 29'h120000e8;
        data[226] = 29'h0b80000f;
        data[227] = 29'h1600f002;
        data[228] = 29'h05ff0001;
        data[229] = 29'h120000e8;
        data[230] = 29'h03ff0001;
        data[231] = 29'h1700f000;
        data[232] = 29'h0f880130;
        data[233] = 29'h15080006;
        data[234] = 29'h0b88fecf;
        data[235] = 29'h15080006;
        data[236] = 29'h18e00009;
        data[237] = 29'h0bee0002;
        data[238] = 29'h120100f0;
        data[239] = 29'h120000ec;
        data[240] = 29'h03ff0001;
        data[241] = 29'h1700f000;
        data[242] = 29'h13100000;
        data[243] = 29'h03000001;
        data[244] = 29'h03110000;
        data[245] = 29'h120100fe;
        data[246] = 29'h0f110100;
        data[247] = 29'h15010006;
        data[248] = 29'h0b1100ff;
        data[249] = 29'h15010006;
        data[250] = 29'h18100009;
        data[251] = 29'h0b110002;
        data[252] = 29'h120100f2;
        data[253] = 29'h120000fa;
        data[254] = 29'h03ff0001;
        data[255] = 29'h1700f000;
        data[256] = 29'h01300000;
        data[257] = 29'h01400000;
        data[258] = 29'h05000000;
        data[259] = 29'h12030105;
        data[260] = 29'h12000107;
        data[261] = 29'h04040000;
        data[262] = 29'h0c333000;
        data[263] = 29'h05110000;
        data[264] = 29'h1203010a;
        data[265] = 29'h1200010c;
        data[266] = 29'h04141000;
        data[267] = 29'h0c333000;
        data[268] = 29'h04a01000;
        data[269] = 29'h10001000;
        data[270] = 29'h10101000;
        data[271] = 29'h10001000;
        data[272] = 29'h05110000;
        data[273] = 29'h12010118;
        data[274] = 29'h0ba10001;
        data[275] = 29'h12010115;
        data[276] = 29'h02440000;
        data[277] = 29'h07000001;
        data[278] = 29'h09110001;
        data[279] = 29'h12000110;
        data[280] = 29'h05330000;
        data[281] = 29'h1201011d;
        data[282] = 29'h04014000;
        data[283] = 29'h03ff0001;
        data[284] = 29'h1700f000;
        data[285] = 29'h0a044000;
        data[286] = 29'h03ff0001;
        data[287] = 29'h1700f000;
        data[288] = 29'h05000003;
        data[289] = 29'h12030123;
        data[290] = 29'h12000120;
        data[291] = 29'h03ff0001;
        data[292] = 29'h1700f000;
        data[293] = 29'h0100000d;
        data[294] = 29'h1600f002;
        data[295] = 29'h05ff0001;
        data[296] = 29'h12000091;
        data[297] = 29'h0100000a;
        data[298] = 29'h1600f002;
        data[299] = 29'h05ff0001;
        data[300] = 29'h12000091;
        data[301] = 29'h01000020;
        data[302] = 29'h1600f002;
        data[303] = 29'h05ff0001;
        data[304] = 29'h12000091;
        data[305] = 29'h0100002d;
        data[306] = 29'h1600f002;
        data[307] = 29'h05ff0001;
        data[308] = 29'h12000091;
        data[309] = 29'h0100002d;
        data[310] = 29'h1600f002;
        data[311] = 29'h05ff0001;
        data[312] = 29'h12000091;
        data[313] = 29'h0100002d;
        data[314] = 29'h1600f002;
        data[315] = 29'h05ff0001;
        data[316] = 29'h12000091;
        data[317] = 29'h01000020;
        data[318] = 29'h1600f002;
        data[319] = 29'h05ff0001;
        data[320] = 29'h12000091;
        data[321] = 29'h01000054;
        data[322] = 29'h1600f002;
        data[323] = 29'h05ff0001;
        data[324] = 29'h12000091;
        data[325] = 29'h01000065;
        data[326] = 29'h1600f002;
        data[327] = 29'h05ff0001;
        data[328] = 29'h12000091;
        data[329] = 29'h01000073;
        data[330] = 29'h1600f002;
        data[331] = 29'h05ff0001;
        data[332] = 29'h12000091;
        data[333] = 29'h01000074;
        data[334] = 29'h1600f002;
        data[335] = 29'h05ff0001;
        data[336] = 29'h12000091;
        data[337] = 29'h01000065;
        data[338] = 29'h1600f002;
        data[339] = 29'h05ff0001;
        data[340] = 29'h12000091;
        data[341] = 29'h01000075;
        data[342] = 29'h1600f002;
        data[343] = 29'h05ff0001;
        data[344] = 29'h12000091;
        data[345] = 29'h01000072;
        data[346] = 29'h1600f002;
        data[347] = 29'h05ff0001;
        data[348] = 29'h12000091;
        data[349] = 29'h01000020;
        data[350] = 29'h1600f002;
        data[351] = 29'h05ff0001;
        data[352] = 29'h12000091;
        data[353] = 29'h01000064;
        data[354] = 29'h1600f002;
        data[355] = 29'h05ff0001;
        data[356] = 29'h12000091;
        data[357] = 29'h01000065;
        data[358] = 29'h1600f002;
        data[359] = 29'h05ff0001;
        data[360] = 29'h12000091;
        data[361] = 29'h01000020;
        data[362] = 29'h1600f002;
        data[363] = 29'h05ff0001;
        data[364] = 29'h12000091;
        data[365] = 29'h01000052;
        data[366] = 29'h1600f002;
        data[367] = 29'h05ff0001;
        data[368] = 29'h12000091;
        data[369] = 29'h01000041;
        data[370] = 29'h1600f002;
        data[371] = 29'h05ff0001;
        data[372] = 29'h12000091;
        data[373] = 29'h0100004d;
        data[374] = 29'h1600f002;
        data[375] = 29'h05ff0001;
        data[376] = 29'h12000091;
        data[377] = 29'h01000020;
        data[378] = 29'h1600f002;
        data[379] = 29'h05ff0001;
        data[380] = 29'h12000091;
        data[381] = 29'h0100002d;
        data[382] = 29'h1600f002;
        data[383] = 29'h05ff0001;
        data[384] = 29'h12000091;
        data[385] = 29'h0100002d;
        data[386] = 29'h1600f002;
        data[387] = 29'h05ff0001;
        data[388] = 29'h12000091;
        data[389] = 29'h0100002d;
        data[390] = 29'h1600f002;
        data[391] = 29'h05ff0001;
        data[392] = 29'h12000091;
        data[393] = 29'h0100000d;
        data[394] = 29'h1600f002;
        data[395] = 29'h05ff0001;
        data[396] = 29'h12000091;
        data[397] = 29'h0100000a;
        data[398] = 29'h1600f002;
        data[399] = 29'h05ff0001;
        data[400] = 29'h12000091;
        data[401] = 29'h0100000d;
        data[402] = 29'h1600f002;
        data[403] = 29'h05ff0001;
        data[404] = 29'h12000091;
        data[405] = 29'h0100000a;
        data[406] = 29'h1600f002;
        data[407] = 29'h05ff0001;
        data[408] = 29'h12000091;
        data[409] = 29'h03ff0001;
        data[410] = 29'h1700f000;
    end
    
    // Lecture synchrone ou asynchrone de la ROM
    always @(*) begin
        DataROM = data[AddrROM];
    end
endmodule
